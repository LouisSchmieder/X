module token

pub struct Position {
pub:
	line_nr u32
	char    u32
	tok     string
}
